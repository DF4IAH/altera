    rom['h 0000] = 32'h EA00_0006;   // addr: 0x0000
    rom['h 0001] = 32'h EAFF_FFFE;   // addr: 0x0004
    rom['h 0002] = 32'h EAFF_FFFE;   // addr: 0x0008
    rom['h 0003] = 32'h EAFF_FFFE;   // addr: 0x000c
    rom['h 0004] = 32'h EAFF_FFFE;   // addr: 0x0010
    rom['h 0005] = 32'h EAFF_FFFE;   // addr: 0x0014
    rom['h 0006] = 32'h EAFF_FFFE;   // addr: 0x0018
    rom['h 0007] = 32'h EAFF_FFFE;   // addr: 0x001c
    rom['h 0008] = 32'h E59F_D004;   // addr: 0x0020
    rom['h 0009] = 32'h EB00_0008;   // addr: 0x0024
    rom['h 0010] = 32'h EAFF_FFFE;   // addr: 0x0028
    rom['h 0011] = 32'h 0000_4000;   // addr: 0x002c
    rom['h 0012] = 32'h E59F_2010;   // addr: 0x0030
    rom['h 0013] = 32'h E592_3000;   // addr: 0x0034
    rom['h 0014] = 32'h E283_1004;   // addr: 0x0038
    rom['h 0015] = 32'h E582_1000;   // addr: 0x003c
    rom['h 0016] = 32'h E583_0000;   // addr: 0x0040
    rom['h 0017] = 32'h E1A0_F00E;   // addr: 0x0044
    rom['h 0018] = 32'h 0000_0098;   // addr: 0x0048
    rom['h 0019] = 32'h E92D_47F0;   // addr: 0x004c
    rom['h 0020] = 32'h E3E0_6002;   // addr: 0x0050
    rom['h 0021] = 32'h E3A0_5009;   // addr: 0x0054
    rom['h 0022] = 32'h E3A0_4000;   // addr: 0x0058
    rom['h 0023] = 32'h E1A0_9005;   // addr: 0x005c
    rom['h 0024] = 32'h E1A0_8004;   // addr: 0x0060
    rom['h 0025] = 32'h E3A0_7003;   // addr: 0x0064
    rom['h 0026] = 32'h E088_8009;   // addr: 0x0068
    rom['h 0027] = 32'h E1A0_0008;   // addr: 0x006c
    rom['h 0028] = 32'h EBFF_FFEE;   // addr: 0x0070
    rom['h 0029] = 32'h E089_9006;   // addr: 0x0074
    rom['h 0030] = 32'h E257_7001;   // addr: 0x0078
    rom['h 0031] = 32'h 1AFF_FFF9;   // addr: 0x007c
    rom['h 0032] = 32'h E084_4085;   // addr: 0x0080
    rom['h 0033] = 32'h E245_5003;   // addr: 0x0084
    rom['h 0034] = 32'h E296_6001;   // addr: 0x0088
    rom['h 0035] = 32'h 1AFF_FFF2;   // addr: 0x008c
    rom['h 0036] = 32'h E1A0_0004;   // addr: 0x0090
    rom['h 0037] = 32'h E8BD_87F0;   // addr: 0x0094
    rom['h 0038] = 32'h 1000_0000;   // addr: 0x0098
